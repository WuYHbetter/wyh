library ieee;
use ieee.std_logic_1164.all;
entity sin2 is
port(clock:in std_logic;
frequence : in std_logic;
dout4:out integer range 0 to 255);
end sin2;
architecture bhv of sin2 is
type mem_type is array(0 to 255) of integer range 0 to 255;
constant mem:mem_type:=(128, 131, 134, 137, 141, 144, 147, 150, 153, 156, 159, 
162, 165, 168, 171, 174, 177, 180, 183, 186, 189, 191, 194, 197, 199, 202, 205,
 207, 209, 212, 214, 217, 219, 221, 223, 225, 227, 229, 231, 233, 235, 236, 238,
  240, 241, 243, 244, 245, 246, 248, 249, 250, 251, 252, 252, 253, 254, 254, 255,
   255, 255, 256, 256, 256, 256, 256, 256, 256, 255, 255, 254, 254, 253, 253, 252,
    251, 250, 249, 248, 247, 246, 245, 243, 242, 240, 239, 237, 236, 234, 232, 230,
     228, 226, 224, 222, 220, 218, 215, 213, 211, 208, 206, 203, 201, 198, 195, 193,
      190, 187, 184, 181, 179, 176, 173, 170, 167, 164, 161, 158, 155, 152, 148, 145,
       142, 139, 136, 133, 130, 126, 123, 120, 117, 114, 111, 108, 104, 101, 98, 95,
        92, 89, 86, 83, 80, 77, 75, 72, 69, 66, 63, 61, 58, 55, 53, 50, 48, 45, 43,
         41, 38, 36, 34, 32, 30, 28, 26, 24, 22, 20, 19, 17, 16, 14, 13, 11, 10,
          9, 8, 7, 6, 5, 4, 3, 3, 2, 2, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 2,
           2, 3, 4, 4, 5, 6, 7, 8, 10, 11, 12, 13, 15, 16, 18, 20, 21, 23, 
           25, 27, 29, 31, 33, 35, 37, 39, 42, 44, 47, 49, 51, 54, 57, 59, 62,
            65, 67, 70, 73, 76, 79, 82, 85, 88, 91, 94, 97, 100, 103, 106, 109,
             112, 115, 119, 122, 125, 128);
signal address:integer range 0 to 255;
begin
 process(clock)
 begin
    if clock'event and clock='1' then
        if (frequence = '0') then
			if address>255 then
				 address<=0;
			else
				 address<=address+1;
				 dout4<=mem(address);
				
			end if;
		else
			if address>=254 then
				 address<=0;
			else
				 address<=address+2;
				 dout4<=mem(address);	
			end if;
		end if;
   end if;
end process;
end bhv;
