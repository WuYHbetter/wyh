library ieee;
use ieee.std_logic_1164.all;
entity fangbo is
port(clock:in std_logic;
frequence : in std_logic;
dout1:out integer range 0 to 255);
end fangbo;
architecture bhv of fangbo is
	type mem_type is array(0 to 255) of integer range 0 to 255;
	constant mem:mem_type:=(50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
	 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
	  50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
	   50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50,
	    50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 50, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 
	    240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240,
	     240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240,
	      240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240,
	       240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240,
	        240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240,
	         240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240, 240,
	          240, 240, 240, 240, 240, 240, 240, 240, 240);
	signal address:integer range 0 to 255;
	
	begin
process(clock)
begin
	if clock'event and clock='1' then
		if (frequence = '0') then
			if address>255 then
				 address<=0;
			else
				 address<=address+1;
				 dout1<=mem(address);
				
			end if;
		else
			if address>=254 then
				 address<=0;
			else
				 address<=address+2;
				 dout1<=mem(address);	
			end if;
		end if;
	end if;
end process;
end bhv;
